
module fpu_wrapper(
  input wire clk,
  input wire [9:0]fpu_in_valid,
  output wire [31:0] fpu_out,
  output wire fpu_out_valid,
  input wire [31:0] fadd_out,
  input wire [31:0] fsub_out,
  input wire [31:0] fmul_out,
  input wire [31:0] fdiv_out,
  input wire [31:0] fsqrt_out,
  input wire [31:0] fabs_out,
  input wire [7:0] fcmp_out,
  input wire [31:0] fftoi_out,
  input wire [31:0] fitof_out,
  output wire fadd_in_valid_a,
  input wire fadd_in_ready_a,
  output wire fadd_in_valid_b,
  input wire fadd_in_ready_b,
  input wire fadd_out_valid,
  output wire fsub_in_valid_a,
  input wire fsub_in_ready_a,
  output wire fsub_in_valid_b,
  input wire fsub_in_ready_b,
  input wire fsub_out_valid,
  output wire fmul_in_valid_a,
  input wire fmul_in_ready_a,
  output wire fmul_in_valid_b,
  input wire fmul_in_ready_b,
  input wire fmul_out_valid,
  output wire fdiv_in_valid_a,
  input wire fdiv_in_ready_a,
  output wire fdiv_in_valid_b,
  input wire fdiv_in_ready_b,
  input wire fdiv_out_valid,
  output wire fsqrt_in_valid_a,
  input wire fsqrt_in_ready_a,
  input wire fsqrt_out_valid,
  output wire fabs_in_valid_a,
  input wire fabs_in_ready_a,
  input wire fabs_out_valid,
  output wire fcmp_in_valid_a,
  input wire fcmp_in_ready_a,
  output wire fcmp_in_valid_b,
  input wire fcmp_in_ready_b,
  output wire fcmp_in_valid_op,
  input wire fcmp_in_ready_op,
  input wire fcmp_out_valid,
  output wire fftoi_in_valid_a,
  input wire fftoi_in_ready_a,
  input wire fftoi_out_valid,
  output wire fitof_in_valid_a,
  input wire fitof_in_ready_a,
  input wire fitof_out_valid
  );

  fpu f1(
    .clk(clk),
    .fpu_in_valid(fpu_in_valid),
    .fpu_out(fpu_out),
    .fpu_out_valid(fpu_out_valid),
    .fadd_out(fadd_out),
    .fsub_out(fsub_out),
    .fmul_out(fmul_out),
    .fdiv_out(fdiv_out),
    .fsqrt_out(fsqrt_out),
    .fabs_out(fabs_out),
    .fcmp_out(fcmp_out),
    .fftoi_out(fftoi_out),
    .fitof_out(fitof_out),
    .fadd_in_valid_a(fadd_in_valid_a),
    .fadd_in_ready_a(fadd_in_ready_a),
    .fadd_in_valid_b(fadd_in_valid_b),
    .fadd_in_ready_b(fadd_in_ready_b),
    .fadd_out_valid(fadd_out_valid),
    .fsub_in_valid_a(fsub_in_valid_a),
    .fsub_in_ready_a(fsub_in_ready_a),
    .fsub_in_valid_b(fsub_in_valid_b),
    .fsub_in_ready_b(fsub_in_ready_b),
    .fsub_out_valid(fsub_out_valid),
    .fmul_in_valid_a(fmul_in_valid_a),
    .fmul_in_ready_a(fmul_in_ready_a),
    .fmul_in_valid_b(fmul_in_valid_b),
    .fmul_in_ready_b(fmul_in_ready_b),
    .fmul_out_valid(fmul_out_valid),
    .fdiv_in_valid_a(fdiv_in_valid_a),
    .fdiv_in_ready_a(fdiv_in_ready_a),
    .fdiv_in_valid_b(fdiv_in_valid_b),
    .fdiv_in_ready_b(fdiv_in_ready_b),
    .fdiv_out_valid(fdiv_out_valid),
    .fsqrt_in_valid_a(fsqrt_in_valid_a),
    .fsqrt_in_ready_a(fsqrt_in_ready_a),
    .fsqrt_out_valid(fsqrt_out_valid),
    .fabs_in_valid_a(fabs_in_valid_a),
    .fabs_in_ready_a(fabs_in_ready_a),
    .fabs_out_valid(fabs_out_valid),
    .fcmp_in_valid_a(fcmp_in_valid_a),
    .fcmp_in_ready_a(fcmp_in_ready_a),
    .fcmp_in_valid_b(fcmp_in_valid_b),
    .fcmp_in_ready_b(fcmp_in_ready_b),
    .fcmp_in_valid_op(fcmp_in_valid_op),
    .fcmp_in_ready_op(fcmp_in_ready_op),
    .fcmp_out_valid(fcmp_out_valid),
    .fftoi_in_valid_a(fftoi_in_valid_a),
    .fftoi_in_ready_a(fftoi_in_ready_a),
    .fftoi_out_valid(fftoi_out_valid),
    .fitof_in_valid_a(fitof_in_valid_a),
    .fitof_in_ready_a(fitof_in_ready_a),
    .fitof_out_valid(fitof_out_valid)
    );

endmodule
