module uart_wrapper (
  input wire clk,
  output wire [3:0] uart_araddr,
  input wire uart_arready,
  output wire uart_arvalid,
  output wire [3:0] uart_awaddr,
  input wire uart_awready,
  output wire uart_awvalid,
  output wire uart_bready,
  input wire [1:0] uart_bresp,
  input wire uart_bvalid,
  input wire [31:0] uart_rdata,
  output wire uart_rready,
  input wire [1:0] uart_rresp,
  input wire uart_rvalid,
  output wire [31:0] uart_wdata,
  input wire uart_wready,
  output wire [3:0] uart_wstrb,
  output wire uart_wvalid,
  input wire [7:0] uart_output,
  input wire uart_outready,
  output wire uart_outvalid,
  output wire [7:0] uart_input,
  input wire uart_inready,
  output wire uart_invalid
  );

  uart u1( clk,
    uart_araddr,
    uart_arready,
    uart_arvalid,
    uart_awaddr,
    uart_awready,
    uart_awvalid,
    uart_bready,
    uart_bresp,
    uart_bvalid,
    uart_rdata,
    uart_rready,
    uart_rresp,
    uart_rvalid,
    uart_wdata,
    uart_wready,
    uart_wstrb,
    uart_wvalid,
    uart_output,
    uart_outready,
    uart_outvalid,
    uart_input,
    uart_inready,
    uart_invalid);

endmodule
